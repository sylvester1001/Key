module display ();




endmodule
