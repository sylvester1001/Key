module mimasuo();




endmodule
